interface XOR_INTF
(
    input logic clk                //signal that will be passed from the top module
);

    logic   A;
    logic   B;
    logic   Y;


endinterface : XOR_INTF
