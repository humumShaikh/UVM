interface ha_intf
(
    input logic clk
);

    logic   A;
    logic   B;
    logic   S;
    logic   C;

endinterface : ha_intf