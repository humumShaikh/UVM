package halfAdder_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "seq_item.sv"
    `include "base_seq.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "environment.sv"

endpackage : halfAdder_pkg