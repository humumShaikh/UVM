module xor_gate
(
    input   logic   A,
    input   logic   B,
    output  logic   Y
);

    assign Y = A ^ B;

endmodule : xor_gate