package xorGate_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "seq_item.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "scoreboard.sv"
    `include "environment.sv"

endpackage : xorGate_pkg