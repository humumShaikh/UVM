interface AND_INTF
(
    input logic clk
);

    logic   A;
    logic   B;
    logic   Y;

endinterface : AND_INTF