interface XOR_INTF
(
    input logic clk
);

    logic   A;
    logic   B;
    logic   Y;

endinterface : XOR_INTF